//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2023 Fall
//   Lab01 Exercise		: Supper MOSFET Calculator
//   Author     		: Lin-Hung Lai (lhlai@ieee.org)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : SMC.v
//   Module Name : SMC
//   Release version : V1.0 (Release Date: 2023-09)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################


module SMC(
  // Input signals
    mode,
    W_0, V_GS_0, V_DS_0,
    W_1, V_GS_1, V_DS_1,
    W_2, V_GS_2, V_DS_2,
    W_3, V_GS_3, V_DS_3,
    W_4, V_GS_4, V_DS_4,
    W_5, V_GS_5, V_DS_5,   
  // Output signals
    out_n
);

//================================================================
//   INPUT AND OUTPUT DECLARATION                         
//================================================================
input [2:0] W_0, V_GS_0, V_DS_0;
input [2:0] W_1, V_GS_1, V_DS_1;
input [2:0] W_2, V_GS_2, V_DS_2;
input [2:0] W_3, V_GS_3, V_DS_3;
input [2:0] W_4, V_GS_4, V_DS_4;
input [2:0] W_5, V_GS_5, V_DS_5;
input [1:0] mode;
output [7:0] out_n;         					// use this if using continuous assignment for out_n  // Ex: assign out_n = XXX;
//output reg [7:0] out_n; 								// use this if using procedure assignment for out_n   // Ex: always@(*) begin out_n = XXX; end

//================================================================
//    Wire & Registers 
//================================================================
// Declare the wire/reg you would use in your circuit
// remember 
// wire for port connection and cont. assignment
// reg for proc. assignment
wire [2:0] W            [0:5];
wire [2:0] V_GS         [0:5];
wire [2:0] V_DS         [0:5];
//  

wire       triode       [0:5];
wire [3:0] id_a         [0:5];
//wire [2:0] id_b         [0:5];
wire [3:0] gm_a         [0:5];
//wire [2:0] gm_b         [0:5];
wire [3:0] mult_a       [0:5];
wire [2:0] mult_b       [0:5];
wire [2:0] mult_c       [0:5]; 
wire [7:0] mult_temp    [0:5];
wire [7:0] mult_result  [0:5];
//sort
wire [7:0] n_0, n_1, n_2, n_3, n_4, n_5;
//
reg [9:0] add_a, add_b, add_c;
//wire [7:0] ave_a, ave_b, ave_c;
//wire [9:0] add_a, add_b, add_c;
wire [9:0] add_result;
wire [9:0] add_temp;


//================================================================
//    Parameter
//================================================================
parameter SIGNAL_NUM = 6;

//================================================================
//    DESIGN
//================================================================

// --------------------------------------------------
// write your design here
// --------------------------------------------------

assign W[0] = W_0;
assign W[1] = W_1;
assign W[2] = W_2;
assign W[3] = W_3;
assign W[4] = W_4;
assign W[5] = W_5;
assign V_GS[0] = V_GS_0;
assign V_GS[1] = V_GS_1;
assign V_GS[2] = V_GS_2;
assign V_GS[3] = V_GS_3;
assign V_GS[4] = V_GS_4;
assign V_GS[5] = V_GS_5;
assign V_DS[0] = V_DS_0;
assign V_DS[1] = V_DS_1;
assign V_DS[2] = V_DS_2;
assign V_DS[3] = V_DS_3;
assign V_DS[4] = V_DS_4;
assign V_DS[5] = V_DS_5;

/*Calculate Id or gm*/

genvar tri_i;
generate
  for(tri_i=0; tri_i < SIGNAL_NUM; tri_i = tri_i+1)begin
    assign triode[tri_i] = (V_GS[tri_i]-1 > V_DS[tri_i]);
  end
endgenerate


genvar id_i;
generate
  for(id_i=0; id_i < SIGNAL_NUM; id_i = id_i+1)begin
    assign id_a[id_i] = (triode[id_i]) ? (2*V_GS[id_i] - 2 - V_DS[id_i]) : (V_GS[id_i] - 1);
  end
endgenerate


genvar gm_i;
generate
  for(gm_i=0; gm_i < SIGNAL_NUM; gm_i = gm_i+1)begin
    assign gm_a[gm_i] = 2;
  end
endgenerate

genvar mult_i;
generate
  for(mult_i=0; mult_i < SIGNAL_NUM; mult_i = mult_i+1)begin
    assign mult_a[mult_i] = (mode[0]) ? id_a[mult_i] : gm_a[mult_i];
    assign mult_b[mult_i] = (triode[mult_i]) ? V_DS[mult_i] : (V_GS[mult_i] - 1);
    assign mult_c[mult_i] = W[mult_i];
  end
endgenerate

generate
  for(mult_i=0; mult_i < SIGNAL_NUM; mult_i = mult_i+1)begin
    assign mult_temp[mult_i] = (mult_a[mult_i] * mult_b[mult_i] * mult_c[mult_i]);
  end
endgenerate

genvar div_i;
generate
  for(div_i=0; div_i < SIGNAL_NUM; div_i = div_i+1)begin
    div_3_in8_out8 u_div_3_in8_out8( .in(mult_temp[div_i]), .out(mult_result[div_i]));
  end
endgenerate

/*
genvar i;
generate
  for(i=0; i < SIGNAL_NUM; i = i+1)begin
    Cal_id_gm u_Cal_id_gm (.mode_0(mode[0]),.w(W[i]),.v_gs(V_GS[i]),.v_ds(V_DS[i]),.mult_result(mult_result[i]));
  end
endgenerate
*/

/*Sort*/
Sort u_sort( .mult_0(mult_result[0]), .mult_1(mult_result[1]), .mult_2(mult_result[2]),
       .mult_3(mult_result[3]), .mult_4(mult_result[4]), .mult_5(mult_result[5]),
       .n_0(n_0), .n_1(n_1), .n_2(n_2), .n_3(n_3), .n_4(n_4), .n_5(n_5)
);
/*Select according to mode*/

always@(*)begin
  case(mode)
    2'b00:begin
      add_a = n_3;
      add_b = n_4;
      add_c = n_5;
    end
    2'b01:begin
      add_a = 3*n_3;
      add_b = 4*n_4;
      add_c = 5*n_5;
    end
    2'b10:begin
      add_a = n_0;
      add_b = n_1;
      add_c = n_2;
    end
    2'b11:begin
      add_a = 3*n_0;
      add_b = 4*n_1;
      add_c = 5*n_2;
    end
  endcase
end

/*
assign ave_a = (mode[1]) ? n_0 : n_3;
assign ave_b = (mode[1]) ? n_1 : n_4;
assign ave_c = (mode[1]) ? n_2 : n_5;
assign add_a = (mode[0]) ? 3*ave_a : ave_a;
assign add_b = (mode[0]) ? 4*ave_b : ave_b;
assign add_c = (mode[0]) ? 5*ave_c : ave_c;
*/

/*Output*/
assign add_temp = (add_a + add_b + add_c);
div_3_in10_out10 u_div_3_in10_out10(.in(add_temp) ,.out(add_result));
assign out_n = (mode[0]) ? add_result[9:2] : add_result[7:0];


endmodule


//================================================================
//   SUB MODULE
//================================================================
/*
module Cal_id_gm(
  // Input signals
  mode_0,
  w,
  v_gs,
  v_ds,
  // Output signals
  mult_result
);
input mode_0;
input [2:0] w, v_gs, v_ds;
output [7:0] mult_result;

wire       triode       ;
wire [3:0] id_a         ;
wire [2:0] id_b         ;
wire [3:0] gm_a         ;
wire [2:0] gm_b         ;
wire [3:0] mult_a       ;
wire [2:0] mult_b       ;
wire [2:0] mult_c       ; 
wire [9:0] mult_temp    ;

assign triode = (v_gs-1 > v_ds);

assign id_a = (triode) ? (2*v_gs - 2 - v_ds) : (v_gs - 1);
assign id_b = (triode) ? v_ds : (v_gs - 1);

assign gm_a = (triode) ? v_ds : (v_gs - 1);
assign gm_b = 2;

assign mult_a = (mode_0) ? id_a : gm_a;
assign mult_b = (mode_0) ? id_b : gm_b;
assign mult_c = w;

assign mult_temp = (mult_a * mult_b * mult_c);

div_3_in10_out8 u_div_3_in10_out8( .in(mult_temp), .out(mult_result));


endmodule
*/
module Sort (
  // Input signals
  mult_0,
  mult_1,
  mult_2,
  mult_3,
  mult_4,
  mult_5,
  // Output signals
  n_0,
  n_1,
  n_2,
  n_3,
  n_4,
  n_5
);
//================================================================
//   INPUT AND OUTPUT DECLARATION                         
//================================================================
input [7:0] mult_0, mult_1, mult_2, mult_3, mult_4, mult_5;
output [7:0] n_0, n_1, n_2, n_3, n_4, n_5;


wire [7:0] L0_0[0:3];
wire [7:0] L0_1[0:2];
wire [7:0] L1_0[0:3];
wire [7:0] L1_1[0:2];
wire [7:0]  L_2[0:3];
wire [7:0]  L_3[0:1]; 

//分成兩個部分各三個比較出大,中,小
//part0
assign L0_0[0] = (mult_0  > mult_1 ) ? mult_0  : mult_1;
assign L0_0[1] = (mult_0  > mult_1 ) ? mult_1  : mult_0;
assign L0_0[2] = (L0_0[1] > mult_2 ) ? L0_0[1] : mult_2;
assign L0_0[3] = (L0_0[1] > mult_2 ) ? mult_2  : L0_0[1];
assign L0_1[0] = (L0_0[0] > L0_0[2]) ? L0_0[0] : L0_0[2];
assign L0_1[1] = (L0_0[0] > L0_0[2]) ? L0_0[2] : L0_0[0];
assign L0_1[2] = L0_0[3];

//part1
assign L1_0[0] = (mult_3  > mult_4 ) ? mult_3  : mult_4;
assign L1_0[1] = (mult_3  > mult_4 ) ? mult_4  : mult_3;
assign L1_0[2] = (L1_0[1] > mult_5 ) ? L1_0[1] : mult_5;
assign L1_0[3] = (L1_0[1] > mult_5 ) ? mult_5  : L1_0[1];
assign L1_1[0] = (L1_0[0] > L1_0[2]) ? L1_0[0] : L1_0[2];
assign L1_1[1] = (L1_0[0] > L1_0[2]) ? L1_0[2] : L1_0[0];
assign L1_1[2] = L1_0[3];

//max & min
assign n_0    = (L0_1[0] > L1_1[0]) ? L0_1[0] : L1_1[0];
assign L_2[0] = (L0_1[0] > L1_1[0]) ? L1_1[0] : L0_1[0];
assign L_2[1] = (L0_1[1] > L1_1[1]) ? L0_1[1] : L1_1[1];
assign L_2[2] = (L0_1[1] > L1_1[1]) ? L1_1[1] : L0_1[1];
assign L_2[3] = (L0_1[2] > L1_1[2]) ? L0_1[2] : L1_1[2];
assign n_5    = (L0_1[2] > L1_1[2]) ? L1_1[2] : L0_1[2];

//second max & second min
assign n_1    = (L_2[0] > L_2[1]) ? L_2[0] : L_2[1];
assign L_3[0] = (L_2[0] > L_2[1]) ? L_2[1] : L_2[0];
assign L_3[1] = (L_2[2] > L_2[3]) ? L_2[2] : L_2[3];
assign n_4    = (L_2[2] > L_2[3]) ? L_2[3] : L_2[2];

//mid
assign n_2    = (L_3[0] > L_3[1]) ? L_3[0] : L_3[1];
assign n_3    = (L_3[0] > L_3[1]) ? L_3[1] : L_3[0];


endmodule

module div_3_in8_out8(
  input  [7:0] in,
  output reg [7:0] out 
);

  always@(*)begin
    case(in)
      8'b00000000:out = 8'd0;
      8'b00000001:out = 8'd0;
      8'b00000010:out = 8'd0;
      8'b00000011:out = 8'd1;
      8'b00000100:out = 8'd1;
      8'b00000101:out = 8'd1;
      8'b00000110:out = 8'd2;
      8'b00000111:out = 8'd2;
      8'b00001000:out = 8'd2;
      8'b00001001:out = 8'd3;
      8'b00001010:out = 8'd3;
      8'b00001011:out = 8'd3;
      8'b00001100:out = 8'd4;
      8'b00001101:out = 8'd4;
      8'b00001110:out = 8'd4;
      8'b00001111:out = 8'd5;
      8'b00010000:out = 8'd5;
      8'b00010001:out = 8'd5;
      8'b00010010:out = 8'd6;
      8'b00010011:out = 8'd6;
      8'b00010100:out = 8'd6;
      8'b00010101:out = 8'd7;
      8'b00010110:out = 8'd7;
      8'b00010111:out = 8'd7;
      8'b00011000:out = 8'd8;
      8'b00011001:out = 8'd8;
      8'b00011010:out = 8'd8;
      8'b00011011:out = 8'd9;
      8'b00011100:out = 8'd9;
      8'b00011101:out = 8'd9;
      8'b00011110:out = 8'd10;
      8'b00011111:out = 8'd10;
      8'b00100000:out = 8'd10;
      8'b00100001:out = 8'd11;
      8'b00100010:out = 8'd11;
      8'b00100011:out = 8'd11;
      8'b00100100:out = 8'd12;
      8'b00100101:out = 8'd12;
      8'b00100110:out = 8'd12;
      8'b00100111:out = 8'd13;
      8'b00101000:out = 8'd13;
      8'b00101001:out = 8'd13;
      8'b00101010:out = 8'd14;
      8'b00101011:out = 8'd14;
      8'b00101100:out = 8'd14;
      8'b00101101:out = 8'd15;
      8'b00101110:out = 8'd15;
      8'b00101111:out = 8'd15;
      8'b00110000:out = 8'd16;
      8'b00110001:out = 8'd16;
      8'b00110010:out = 8'd16;
      8'b00110011:out = 8'd17;
      8'b00110100:out = 8'd17;
      8'b00110101:out = 8'd17;
      8'b00110110:out = 8'd18;
      8'b00110111:out = 8'd18;
      8'b00111000:out = 8'd18;
      8'b00111001:out = 8'd19;
      8'b00111010:out = 8'd19;
      8'b00111011:out = 8'd19;
      8'b00111100:out = 8'd20;
      8'b00111101:out = 8'd20;
      8'b00111110:out = 8'd20;
      8'b00111111:out = 8'd21;
      8'b01000000:out = 8'd21;
      8'b01000001:out = 8'd21;
      8'b01000010:out = 8'd22;
      8'b01000011:out = 8'd22;
      8'b01000100:out = 8'd22;
      8'b01000101:out = 8'd23;
      8'b01000110:out = 8'd23;
      8'b01000111:out = 8'd23;
      8'b01001000:out = 8'd24;
      8'b01001001:out = 8'd24;
      8'b01001010:out = 8'd24;
      8'b01001011:out = 8'd25;
      8'b01001100:out = 8'd25;
      8'b01001101:out = 8'd25;
      8'b01001110:out = 8'd26;
      8'b01001111:out = 8'd26;
      8'b01010000:out = 8'd26;
      8'b01010001:out = 8'd27;
      8'b01010010:out = 8'd27;
      8'b01010011:out = 8'd27;
      8'b01010100:out = 8'd28;
      8'b01010101:out = 8'd28;
      8'b01010110:out = 8'd28;
      8'b01010111:out = 8'd29;
      8'b01011000:out = 8'd29;
      8'b01011001:out = 8'd29;
      8'b01011010:out = 8'd30;
      8'b01011011:out = 8'd30;
      8'b01011100:out = 8'd30;
      8'b01011101:out = 8'd31;
      8'b01011110:out = 8'd31;
      8'b01011111:out = 8'd31;
      8'b01100000:out = 8'd32;
      8'b01100001:out = 8'd32;
      8'b01100010:out = 8'd32;
      8'b01100011:out = 8'd33;
      8'b01100100:out = 8'd33;
      8'b01100101:out = 8'd33;
      8'b01100110:out = 8'd34;
      8'b01100111:out = 8'd34;
      8'b01101000:out = 8'd34;
      8'b01101001:out = 8'd35;
      8'b01101010:out = 8'd35;
      8'b01101011:out = 8'd35;
      8'b01101100:out = 8'd36;
      8'b01101101:out = 8'd36;
      8'b01101110:out = 8'd36;
      8'b01101111:out = 8'd37;
      8'b01110000:out = 8'd37;
      8'b01110001:out = 8'd37;
      8'b01110010:out = 8'd38;
      8'b01110011:out = 8'd38;
      8'b01110100:out = 8'd38;
      8'b01110101:out = 8'd39;
      8'b01110110:out = 8'd39;
      8'b01110111:out = 8'd39;
      8'b01111000:out = 8'd40;
      8'b01111001:out = 8'd40;
      8'b01111010:out = 8'd40;
      8'b01111011:out = 8'd41;
      8'b01111100:out = 8'd41;
      8'b01111101:out = 8'd41;
      8'b01111110:out = 8'd42;
      8'b01111111:out = 8'd42;
      8'b10000000:out = 8'd42;
      8'b10000001:out = 8'd43;
      8'b10000010:out = 8'd43;
      8'b10000011:out = 8'd43;
      8'b10000100:out = 8'd44;
      8'b10000101:out = 8'd44;
      8'b10000110:out = 8'd44;
      8'b10000111:out = 8'd45;
      8'b10001000:out = 8'd45;
      8'b10001001:out = 8'd45;
      8'b10001010:out = 8'd46;
      8'b10001011:out = 8'd46;
      8'b10001100:out = 8'd46;
      8'b10001101:out = 8'd47;
      8'b10001110:out = 8'd47;
      8'b10001111:out = 8'd47;
      8'b10010000:out = 8'd48;
      8'b10010001:out = 8'd48;
      8'b10010010:out = 8'd48;
      8'b10010011:out = 8'd49;
      8'b10010100:out = 8'd49;
      8'b10010101:out = 8'd49;
      8'b10010110:out = 8'd50;
      8'b10010111:out = 8'd50;
      8'b10011000:out = 8'd50;
      8'b10011001:out = 8'd51;
      8'b10011010:out = 8'd51;
      8'b10011011:out = 8'd51;
      8'b10011100:out = 8'd52;
      8'b10011101:out = 8'd52;
      8'b10011110:out = 8'd52;
      8'b10011111:out = 8'd53;
      8'b10100000:out = 8'd53;
      8'b10100001:out = 8'd53;
      8'b10100010:out = 8'd54;
      8'b10100011:out = 8'd54;
      8'b10100100:out = 8'd54;
      8'b10100101:out = 8'd55;
      8'b10100110:out = 8'd55;
      8'b10100111:out = 8'd55;
      8'b10101000:out = 8'd56;
      8'b10101001:out = 8'd56;
      8'b10101010:out = 8'd56;
      8'b10101011:out = 8'd57;
      8'b10101100:out = 8'd57;
      8'b10101101:out = 8'd57;
      8'b10101110:out = 8'd58;
      8'b10101111:out = 8'd58;
      8'b10110000:out = 8'd58;
      8'b10110001:out = 8'd59;
      8'b10110010:out = 8'd59;
      8'b10110011:out = 8'd59;
      8'b10110100:out = 8'd60;
      8'b10110101:out = 8'd60;
      8'b10110110:out = 8'd60;
      8'b10110111:out = 8'd61;
      8'b10111000:out = 8'd61;
      8'b10111001:out = 8'd61;
      8'b10111010:out = 8'd62;
      8'b10111011:out = 8'd62;
      8'b10111100:out = 8'd62;
      8'b10111101:out = 8'd63;
      8'b10111110:out = 8'd63;
      8'b10111111:out = 8'd63;
      8'b11000000:out = 8'd64;
      8'b11000001:out = 8'd64;
      8'b11000010:out = 8'd64;
      8'b11000011:out = 8'd65;
      8'b11000100:out = 8'd65;
      8'b11000101:out = 8'd65;
      8'b11000110:out = 8'd66;
      8'b11000111:out = 8'd66;
      8'b11001000:out = 8'd66;
      8'b11001001:out = 8'd67;
      8'b11001010:out = 8'd67;
      8'b11001011:out = 8'd67;
      8'b11001100:out = 8'd68;
      8'b11001101:out = 8'd68;
      8'b11001110:out = 8'd68;
      8'b11001111:out = 8'd69;
      8'b11010000:out = 8'd69;
      8'b11010001:out = 8'd69;
      8'b11010010:out = 8'd70;
      8'b11010011:out = 8'd70;
      8'b11010100:out = 8'd70;
      8'b11010101:out = 8'd71;
      8'b11010110:out = 8'd71;
      8'b11010111:out = 8'd71;
      8'b11011000:out = 8'd72;
      8'b11011001:out = 8'd72;
      8'b11011010:out = 8'd72;
      8'b11011011:out = 8'd73;
      8'b11011100:out = 8'd73;
      8'b11011101:out = 8'd73;
      8'b11011110:out = 8'd74;
      8'b11011111:out = 8'd74;
      8'b11100000:out = 8'd74;
      8'b11100001:out = 8'd75;
      8'b11100010:out = 8'd75;
      8'b11100011:out = 8'd75;
      8'b11100100:out = 8'd76;
      8'b11100101:out = 8'd76;
      8'b11100110:out = 8'd76;
      8'b11100111:out = 8'd77;
      8'b11101000:out = 8'd77;
      8'b11101001:out = 8'd77;
      8'b11101010:out = 8'd78;
      8'b11101011:out = 8'd78;
      8'b11101100:out = 8'd78;
      8'b11101101:out = 8'd79;
      8'b11101110:out = 8'd79;
      8'b11101111:out = 8'd79;
      8'b11110000:out = 8'd80;
      8'b11110001:out = 8'd80;
      8'b11110010:out = 8'd80;
      8'b11110011:out = 8'd81;
      8'b11110100:out = 8'd81;
      8'b11110101:out = 8'd81;
      8'b11110110:out = 8'd82;
      8'b11110111:out = 8'd82;
      8'b11111000:out = 8'd82;
      8'b11111001:out = 8'd83;
      8'b11111010:out = 8'd83;
      8'b11111011:out = 8'd83;
      8'b11111100:out = 8'd84;
      8'b11111101:out = 8'd84;
      8'b11111110:out = 8'd84;
      8'b11111111:out = 8'd85;
    endcase
  end
endmodule

module div_3_in10_out10(
  input  [9:0] in,
  output reg [9:0] out 
);

  always@(*)begin
    case(in)
      10'b0000000000:out = 10'd0;
      10'b0000000001:out = 10'd0;
      10'b0000000010:out = 10'd0;
      10'b0000000011:out = 10'd1;
      10'b0000000100:out = 10'd1;
      10'b0000000101:out = 10'd1;
      10'b0000000110:out = 10'd2;
      10'b0000000111:out = 10'd2;
      10'b0000001000:out = 10'd2;
      10'b0000001001:out = 10'd3;
      10'b0000001010:out = 10'd3;
      10'b0000001011:out = 10'd3;
      10'b0000001100:out = 10'd4;
      10'b0000001101:out = 10'd4;
      10'b0000001110:out = 10'd4;
      10'b0000001111:out = 10'd5;
      10'b0000010000:out = 10'd5;
      10'b0000010001:out = 10'd5;
      10'b0000010010:out = 10'd6;
      10'b0000010011:out = 10'd6;
      10'b0000010100:out = 10'd6;
      10'b0000010101:out = 10'd7;
      10'b0000010110:out = 10'd7;
      10'b0000010111:out = 10'd7;
      10'b0000011000:out = 10'd8;
      10'b0000011001:out = 10'd8;
      10'b0000011010:out = 10'd8;
      10'b0000011011:out = 10'd9;
      10'b0000011100:out = 10'd9;
      10'b0000011101:out = 10'd9;
      10'b0000011110:out = 10'd10;
      10'b0000011111:out = 10'd10;
      10'b0000100000:out = 10'd10;
      10'b0000100001:out = 10'd11;
      10'b0000100010:out = 10'd11;
      10'b0000100011:out = 10'd11;
      10'b0000100100:out = 10'd12;
      10'b0000100101:out = 10'd12;
      10'b0000100110:out = 10'd12;
      10'b0000100111:out = 10'd13;
      10'b0000101000:out = 10'd13;
      10'b0000101001:out = 10'd13;
      10'b0000101010:out = 10'd14;
      10'b0000101011:out = 10'd14;
      10'b0000101100:out = 10'd14;
      10'b0000101101:out = 10'd15;
      10'b0000101110:out = 10'd15;
      10'b0000101111:out = 10'd15;
      10'b0000110000:out = 10'd16;
      10'b0000110001:out = 10'd16;
      10'b0000110010:out = 10'd16;
      10'b0000110011:out = 10'd17;
      10'b0000110100:out = 10'd17;
      10'b0000110101:out = 10'd17;
      10'b0000110110:out = 10'd18;
      10'b0000110111:out = 10'd18;
      10'b0000111000:out = 10'd18;
      10'b0000111001:out = 10'd19;
      10'b0000111010:out = 10'd19;
      10'b0000111011:out = 10'd19;
      10'b0000111100:out = 10'd20;
      10'b0000111101:out = 10'd20;
      10'b0000111110:out = 10'd20;
      10'b0000111111:out = 10'd21;
      10'b0001000000:out = 10'd21;
      10'b0001000001:out = 10'd21;
      10'b0001000010:out = 10'd22;
      10'b0001000011:out = 10'd22;
      10'b0001000100:out = 10'd22;
      10'b0001000101:out = 10'd23;
      10'b0001000110:out = 10'd23;
      10'b0001000111:out = 10'd23;
      10'b0001001000:out = 10'd24;
      10'b0001001001:out = 10'd24;
      10'b0001001010:out = 10'd24;
      10'b0001001011:out = 10'd25;
      10'b0001001100:out = 10'd25;
      10'b0001001101:out = 10'd25;
      10'b0001001110:out = 10'd26;
      10'b0001001111:out = 10'd26;
      10'b0001010000:out = 10'd26;
      10'b0001010001:out = 10'd27;
      10'b0001010010:out = 10'd27;
      10'b0001010011:out = 10'd27;
      10'b0001010100:out = 10'd28;
      10'b0001010101:out = 10'd28;
      10'b0001010110:out = 10'd28;
      10'b0001010111:out = 10'd29;
      10'b0001011000:out = 10'd29;
      10'b0001011001:out = 10'd29;
      10'b0001011010:out = 10'd30;
      10'b0001011011:out = 10'd30;
      10'b0001011100:out = 10'd30;
      10'b0001011101:out = 10'd31;
      10'b0001011110:out = 10'd31;
      10'b0001011111:out = 10'd31;
      10'b0001100000:out = 10'd32;
      10'b0001100001:out = 10'd32;
      10'b0001100010:out = 10'd32;
      10'b0001100011:out = 10'd33;
      10'b0001100100:out = 10'd33;
      10'b0001100101:out = 10'd33;
      10'b0001100110:out = 10'd34;
      10'b0001100111:out = 10'd34;
      10'b0001101000:out = 10'd34;
      10'b0001101001:out = 10'd35;
      10'b0001101010:out = 10'd35;
      10'b0001101011:out = 10'd35;
      10'b0001101100:out = 10'd36;
      10'b0001101101:out = 10'd36;
      10'b0001101110:out = 10'd36;
      10'b0001101111:out = 10'd37;
      10'b0001110000:out = 10'd37;
      10'b0001110001:out = 10'd37;
      10'b0001110010:out = 10'd38;
      10'b0001110011:out = 10'd38;
      10'b0001110100:out = 10'd38;
      10'b0001110101:out = 10'd39;
      10'b0001110110:out = 10'd39;
      10'b0001110111:out = 10'd39;
      10'b0001111000:out = 10'd40;
      10'b0001111001:out = 10'd40;
      10'b0001111010:out = 10'd40;
      10'b0001111011:out = 10'd41;
      10'b0001111100:out = 10'd41;
      10'b0001111101:out = 10'd41;
      10'b0001111110:out = 10'd42;
      10'b0001111111:out = 10'd42;
      10'b0010000000:out = 10'd42;
      10'b0010000001:out = 10'd43;
      10'b0010000010:out = 10'd43;
      10'b0010000011:out = 10'd43;
      10'b0010000100:out = 10'd44;
      10'b0010000101:out = 10'd44;
      10'b0010000110:out = 10'd44;
      10'b0010000111:out = 10'd45;
      10'b0010001000:out = 10'd45;
      10'b0010001001:out = 10'd45;
      10'b0010001010:out = 10'd46;
      10'b0010001011:out = 10'd46;
      10'b0010001100:out = 10'd46;
      10'b0010001101:out = 10'd47;
      10'b0010001110:out = 10'd47;
      10'b0010001111:out = 10'd47;
      10'b0010010000:out = 10'd48;
      10'b0010010001:out = 10'd48;
      10'b0010010010:out = 10'd48;
      10'b0010010011:out = 10'd49;
      10'b0010010100:out = 10'd49;
      10'b0010010101:out = 10'd49;
      10'b0010010110:out = 10'd50;
      10'b0010010111:out = 10'd50;
      10'b0010011000:out = 10'd50;
      10'b0010011001:out = 10'd51;
      10'b0010011010:out = 10'd51;
      10'b0010011011:out = 10'd51;
      10'b0010011100:out = 10'd52;
      10'b0010011101:out = 10'd52;
      10'b0010011110:out = 10'd52;
      10'b0010011111:out = 10'd53;
      10'b0010100000:out = 10'd53;
      10'b0010100001:out = 10'd53;
      10'b0010100010:out = 10'd54;
      10'b0010100011:out = 10'd54;
      10'b0010100100:out = 10'd54;
      10'b0010100101:out = 10'd55;
      10'b0010100110:out = 10'd55;
      10'b0010100111:out = 10'd55;
      10'b0010101000:out = 10'd56;
      10'b0010101001:out = 10'd56;
      10'b0010101010:out = 10'd56;
      10'b0010101011:out = 10'd57;
      10'b0010101100:out = 10'd57;
      10'b0010101101:out = 10'd57;
      10'b0010101110:out = 10'd58;
      10'b0010101111:out = 10'd58;
      10'b0010110000:out = 10'd58;
      10'b0010110001:out = 10'd59;
      10'b0010110010:out = 10'd59;
      10'b0010110011:out = 10'd59;
      10'b0010110100:out = 10'd60;
      10'b0010110101:out = 10'd60;
      10'b0010110110:out = 10'd60;
      10'b0010110111:out = 10'd61;
      10'b0010111000:out = 10'd61;
      10'b0010111001:out = 10'd61;
      10'b0010111010:out = 10'd62;
      10'b0010111011:out = 10'd62;
      10'b0010111100:out = 10'd62;
      10'b0010111101:out = 10'd63;
      10'b0010111110:out = 10'd63;
      10'b0010111111:out = 10'd63;
      10'b0011000000:out = 10'd64;
      10'b0011000001:out = 10'd64;
      10'b0011000010:out = 10'd64;
      10'b0011000011:out = 10'd65;
      10'b0011000100:out = 10'd65;
      10'b0011000101:out = 10'd65;
      10'b0011000110:out = 10'd66;
      10'b0011000111:out = 10'd66;
      10'b0011001000:out = 10'd66;
      10'b0011001001:out = 10'd67;
      10'b0011001010:out = 10'd67;
      10'b0011001011:out = 10'd67;
      10'b0011001100:out = 10'd68;
      10'b0011001101:out = 10'd68;
      10'b0011001110:out = 10'd68;
      10'b0011001111:out = 10'd69;
      10'b0011010000:out = 10'd69;
      10'b0011010001:out = 10'd69;
      10'b0011010010:out = 10'd70;
      10'b0011010011:out = 10'd70;
      10'b0011010100:out = 10'd70;
      10'b0011010101:out = 10'd71;
      10'b0011010110:out = 10'd71;
      10'b0011010111:out = 10'd71;
      10'b0011011000:out = 10'd72;
      10'b0011011001:out = 10'd72;
      10'b0011011010:out = 10'd72;
      10'b0011011011:out = 10'd73;
      10'b0011011100:out = 10'd73;
      10'b0011011101:out = 10'd73;
      10'b0011011110:out = 10'd74;
      10'b0011011111:out = 10'd74;
      10'b0011100000:out = 10'd74;
      10'b0011100001:out = 10'd75;
      10'b0011100010:out = 10'd75;
      10'b0011100011:out = 10'd75;
      10'b0011100100:out = 10'd76;
      10'b0011100101:out = 10'd76;
      10'b0011100110:out = 10'd76;
      10'b0011100111:out = 10'd77;
      10'b0011101000:out = 10'd77;
      10'b0011101001:out = 10'd77;
      10'b0011101010:out = 10'd78;
      10'b0011101011:out = 10'd78;
      10'b0011101100:out = 10'd78;
      10'b0011101101:out = 10'd79;
      10'b0011101110:out = 10'd79;
      10'b0011101111:out = 10'd79;
      10'b0011110000:out = 10'd80;
      10'b0011110001:out = 10'd80;
      10'b0011110010:out = 10'd80;
      10'b0011110011:out = 10'd81;
      10'b0011110100:out = 10'd81;
      10'b0011110101:out = 10'd81;
      10'b0011110110:out = 10'd82;
      10'b0011110111:out = 10'd82;
      10'b0011111000:out = 10'd82;
      10'b0011111001:out = 10'd83;
      10'b0011111010:out = 10'd83;
      10'b0011111011:out = 10'd83;
      10'b0011111100:out = 10'd84;
      10'b0011111101:out = 10'd84;
      10'b0011111110:out = 10'd84;
      10'b0011111111:out = 10'd85;
      10'b0100000000:out = 10'd85;
      10'b0100000001:out = 10'd85;
      10'b0100000010:out = 10'd86;
      10'b0100000011:out = 10'd86;
      10'b0100000100:out = 10'd86;
      10'b0100000101:out = 10'd87;
      10'b0100000110:out = 10'd87;
      10'b0100000111:out = 10'd87;
      10'b0100001000:out = 10'd88;
      10'b0100001001:out = 10'd88;
      10'b0100001010:out = 10'd88;
      10'b0100001011:out = 10'd89;
      10'b0100001100:out = 10'd89;
      10'b0100001101:out = 10'd89;
      10'b0100001110:out = 10'd90;
      10'b0100001111:out = 10'd90;
      10'b0100010000:out = 10'd90;
      10'b0100010001:out = 10'd91;
      10'b0100010010:out = 10'd91;
      10'b0100010011:out = 10'd91;
      10'b0100010100:out = 10'd92;
      10'b0100010101:out = 10'd92;
      10'b0100010110:out = 10'd92;
      10'b0100010111:out = 10'd93;
      10'b0100011000:out = 10'd93;
      10'b0100011001:out = 10'd93;
      10'b0100011010:out = 10'd94;
      10'b0100011011:out = 10'd94;
      10'b0100011100:out = 10'd94;
      10'b0100011101:out = 10'd95;
      10'b0100011110:out = 10'd95;
      10'b0100011111:out = 10'd95;
      10'b0100100000:out = 10'd96;
      10'b0100100001:out = 10'd96;
      10'b0100100010:out = 10'd96;
      10'b0100100011:out = 10'd97;
      10'b0100100100:out = 10'd97;
      10'b0100100101:out = 10'd97;
      10'b0100100110:out = 10'd98;
      10'b0100100111:out = 10'd98;
      10'b0100101000:out = 10'd98;
      10'b0100101001:out = 10'd99;
      10'b0100101010:out = 10'd99;
      10'b0100101011:out = 10'd99;
      10'b0100101100:out = 10'd100;
      10'b0100101101:out = 10'd100;
      10'b0100101110:out = 10'd100;
      10'b0100101111:out = 10'd101;
      10'b0100110000:out = 10'd101;
      10'b0100110001:out = 10'd101;
      10'b0100110010:out = 10'd102;
      10'b0100110011:out = 10'd102;
      10'b0100110100:out = 10'd102;
      10'b0100110101:out = 10'd103;
      10'b0100110110:out = 10'd103;
      10'b0100110111:out = 10'd103;
      10'b0100111000:out = 10'd104;
      10'b0100111001:out = 10'd104;
      10'b0100111010:out = 10'd104;
      10'b0100111011:out = 10'd105;
      10'b0100111100:out = 10'd105;
      10'b0100111101:out = 10'd105;
      10'b0100111110:out = 10'd106;
      10'b0100111111:out = 10'd106;
      10'b0101000000:out = 10'd106;
      10'b0101000001:out = 10'd107;
      10'b0101000010:out = 10'd107;
      10'b0101000011:out = 10'd107;
      10'b0101000100:out = 10'd108;
      10'b0101000101:out = 10'd108;
      10'b0101000110:out = 10'd108;
      10'b0101000111:out = 10'd109;
      10'b0101001000:out = 10'd109;
      10'b0101001001:out = 10'd109;
      10'b0101001010:out = 10'd110;
      10'b0101001011:out = 10'd110;
      10'b0101001100:out = 10'd110;
      10'b0101001101:out = 10'd111;
      10'b0101001110:out = 10'd111;
      10'b0101001111:out = 10'd111;
      10'b0101010000:out = 10'd112;
      10'b0101010001:out = 10'd112;
      10'b0101010010:out = 10'd112;
      10'b0101010011:out = 10'd113;
      10'b0101010100:out = 10'd113;
      10'b0101010101:out = 10'd113;
      10'b0101010110:out = 10'd114;
      10'b0101010111:out = 10'd114;
      10'b0101011000:out = 10'd114;
      10'b0101011001:out = 10'd115;
      10'b0101011010:out = 10'd115;
      10'b0101011011:out = 10'd115;
      10'b0101011100:out = 10'd116;
      10'b0101011101:out = 10'd116;
      10'b0101011110:out = 10'd116;
      10'b0101011111:out = 10'd117;
      10'b0101100000:out = 10'd117;
      10'b0101100001:out = 10'd117;
      10'b0101100010:out = 10'd118;
      10'b0101100011:out = 10'd118;
      10'b0101100100:out = 10'd118;
      10'b0101100101:out = 10'd119;
      10'b0101100110:out = 10'd119;
      10'b0101100111:out = 10'd119;
      10'b0101101000:out = 10'd120;
      10'b0101101001:out = 10'd120;
      10'b0101101010:out = 10'd120;
      10'b0101101011:out = 10'd121;
      10'b0101101100:out = 10'd121;
      10'b0101101101:out = 10'd121;
      10'b0101101110:out = 10'd122;
      10'b0101101111:out = 10'd122;
      10'b0101110000:out = 10'd122;
      10'b0101110001:out = 10'd123;
      10'b0101110010:out = 10'd123;
      10'b0101110011:out = 10'd123;
      10'b0101110100:out = 10'd124;
      10'b0101110101:out = 10'd124;
      10'b0101110110:out = 10'd124;
      10'b0101110111:out = 10'd125;
      10'b0101111000:out = 10'd125;
      10'b0101111001:out = 10'd125;
      10'b0101111010:out = 10'd126;
      10'b0101111011:out = 10'd126;
      10'b0101111100:out = 10'd126;
      10'b0101111101:out = 10'd127;
      10'b0101111110:out = 10'd127;
      10'b0101111111:out = 10'd127;
      10'b0110000000:out = 10'd128;
      10'b0110000001:out = 10'd128;
      10'b0110000010:out = 10'd128;
      10'b0110000011:out = 10'd129;
      10'b0110000100:out = 10'd129;
      10'b0110000101:out = 10'd129;
      10'b0110000110:out = 10'd130;
      10'b0110000111:out = 10'd130;
      10'b0110001000:out = 10'd130;
      10'b0110001001:out = 10'd131;
      10'b0110001010:out = 10'd131;
      10'b0110001011:out = 10'd131;
      10'b0110001100:out = 10'd132;
      10'b0110001101:out = 10'd132;
      10'b0110001110:out = 10'd132;
      10'b0110001111:out = 10'd133;
      10'b0110010000:out = 10'd133;
      10'b0110010001:out = 10'd133;
      10'b0110010010:out = 10'd134;
      10'b0110010011:out = 10'd134;
      10'b0110010100:out = 10'd134;
      10'b0110010101:out = 10'd135;
      10'b0110010110:out = 10'd135;
      10'b0110010111:out = 10'd135;
      10'b0110011000:out = 10'd136;
      10'b0110011001:out = 10'd136;
      10'b0110011010:out = 10'd136;
      10'b0110011011:out = 10'd137;
      10'b0110011100:out = 10'd137;
      10'b0110011101:out = 10'd137;
      10'b0110011110:out = 10'd138;
      10'b0110011111:out = 10'd138;
      10'b0110100000:out = 10'd138;
      10'b0110100001:out = 10'd139;
      10'b0110100010:out = 10'd139;
      10'b0110100011:out = 10'd139;
      10'b0110100100:out = 10'd140;
      10'b0110100101:out = 10'd140;
      10'b0110100110:out = 10'd140;
      10'b0110100111:out = 10'd141;
      10'b0110101000:out = 10'd141;
      10'b0110101001:out = 10'd141;
      10'b0110101010:out = 10'd142;
      10'b0110101011:out = 10'd142;
      10'b0110101100:out = 10'd142;
      10'b0110101101:out = 10'd143;
      10'b0110101110:out = 10'd143;
      10'b0110101111:out = 10'd143;
      10'b0110110000:out = 10'd144;
      10'b0110110001:out = 10'd144;
      10'b0110110010:out = 10'd144;
      10'b0110110011:out = 10'd145;
      10'b0110110100:out = 10'd145;
      10'b0110110101:out = 10'd145;
      10'b0110110110:out = 10'd146;
      10'b0110110111:out = 10'd146;
      10'b0110111000:out = 10'd146;
      10'b0110111001:out = 10'd147;
      10'b0110111010:out = 10'd147;
      10'b0110111011:out = 10'd147;
      10'b0110111100:out = 10'd148;
      10'b0110111101:out = 10'd148;
      10'b0110111110:out = 10'd148;
      10'b0110111111:out = 10'd149;
      10'b0111000000:out = 10'd149;
      10'b0111000001:out = 10'd149;
      10'b0111000010:out = 10'd150;
      10'b0111000011:out = 10'd150;
      10'b0111000100:out = 10'd150;
      10'b0111000101:out = 10'd151;
      10'b0111000110:out = 10'd151;
      10'b0111000111:out = 10'd151;
      10'b0111001000:out = 10'd152;
      10'b0111001001:out = 10'd152;
      10'b0111001010:out = 10'd152;
      10'b0111001011:out = 10'd153;
      10'b0111001100:out = 10'd153;
      10'b0111001101:out = 10'd153;
      10'b0111001110:out = 10'd154;
      10'b0111001111:out = 10'd154;
      10'b0111010000:out = 10'd154;
      10'b0111010001:out = 10'd155;
      10'b0111010010:out = 10'd155;
      10'b0111010011:out = 10'd155;
      10'b0111010100:out = 10'd156;
      10'b0111010101:out = 10'd156;
      10'b0111010110:out = 10'd156;
      10'b0111010111:out = 10'd157;
      10'b0111011000:out = 10'd157;
      10'b0111011001:out = 10'd157;
      10'b0111011010:out = 10'd158;
      10'b0111011011:out = 10'd158;
      10'b0111011100:out = 10'd158;
      10'b0111011101:out = 10'd159;
      10'b0111011110:out = 10'd159;
      10'b0111011111:out = 10'd159;
      10'b0111100000:out = 10'd160;
      10'b0111100001:out = 10'd160;
      10'b0111100010:out = 10'd160;
      10'b0111100011:out = 10'd161;
      10'b0111100100:out = 10'd161;
      10'b0111100101:out = 10'd161;
      10'b0111100110:out = 10'd162;
      10'b0111100111:out = 10'd162;
      10'b0111101000:out = 10'd162;
      10'b0111101001:out = 10'd163;
      10'b0111101010:out = 10'd163;
      10'b0111101011:out = 10'd163;
      10'b0111101100:out = 10'd164;
      10'b0111101101:out = 10'd164;
      10'b0111101110:out = 10'd164;
      10'b0111101111:out = 10'd165;
      10'b0111110000:out = 10'd165;
      10'b0111110001:out = 10'd165;
      10'b0111110010:out = 10'd166;
      10'b0111110011:out = 10'd166;
      10'b0111110100:out = 10'd166;
      10'b0111110101:out = 10'd167;
      10'b0111110110:out = 10'd167;
      10'b0111110111:out = 10'd167;
      10'b0111111000:out = 10'd168;
      10'b0111111001:out = 10'd168;
      10'b0111111010:out = 10'd168;
      10'b0111111011:out = 10'd169;
      10'b0111111100:out = 10'd169;
      10'b0111111101:out = 10'd169;
      10'b0111111110:out = 10'd170;
      10'b0111111111:out = 10'd170;
      10'b1000000000:out = 10'd170;
      10'b1000000001:out = 10'd171;
      10'b1000000010:out = 10'd171;
      10'b1000000011:out = 10'd171;
      10'b1000000100:out = 10'd172;
      10'b1000000101:out = 10'd172;
      10'b1000000110:out = 10'd172;
      10'b1000000111:out = 10'd173;
      10'b1000001000:out = 10'd173;
      10'b1000001001:out = 10'd173;
      10'b1000001010:out = 10'd174;
      10'b1000001011:out = 10'd174;
      10'b1000001100:out = 10'd174;
      10'b1000001101:out = 10'd175;
      10'b1000001110:out = 10'd175;
      10'b1000001111:out = 10'd175;
      10'b1000010000:out = 10'd176;
      10'b1000010001:out = 10'd176;
      10'b1000010010:out = 10'd176;
      10'b1000010011:out = 10'd177;
      10'b1000010100:out = 10'd177;
      10'b1000010101:out = 10'd177;
      10'b1000010110:out = 10'd178;
      10'b1000010111:out = 10'd178;
      10'b1000011000:out = 10'd178;
      10'b1000011001:out = 10'd179;
      10'b1000011010:out = 10'd179;
      10'b1000011011:out = 10'd179;
      10'b1000011100:out = 10'd180;
      10'b1000011101:out = 10'd180;
      10'b1000011110:out = 10'd180;
      10'b1000011111:out = 10'd181;
      10'b1000100000:out = 10'd181;
      10'b1000100001:out = 10'd181;
      10'b1000100010:out = 10'd182;
      10'b1000100011:out = 10'd182;
      10'b1000100100:out = 10'd182;
      10'b1000100101:out = 10'd183;
      10'b1000100110:out = 10'd183;
      10'b1000100111:out = 10'd183;
      10'b1000101000:out = 10'd184;
      10'b1000101001:out = 10'd184;
      10'b1000101010:out = 10'd184;
      10'b1000101011:out = 10'd185;
      10'b1000101100:out = 10'd185;
      10'b1000101101:out = 10'd185;
      10'b1000101110:out = 10'd186;
      10'b1000101111:out = 10'd186;
      10'b1000110000:out = 10'd186;
      10'b1000110001:out = 10'd187;
      10'b1000110010:out = 10'd187;
      10'b1000110011:out = 10'd187;
      10'b1000110100:out = 10'd188;
      10'b1000110101:out = 10'd188;
      10'b1000110110:out = 10'd188;
      10'b1000110111:out = 10'd189;
      10'b1000111000:out = 10'd189;
      10'b1000111001:out = 10'd189;
      10'b1000111010:out = 10'd190;
      10'b1000111011:out = 10'd190;
      10'b1000111100:out = 10'd190;
      10'b1000111101:out = 10'd191;
      10'b1000111110:out = 10'd191;
      10'b1000111111:out = 10'd191;
      10'b1001000000:out = 10'd192;
      10'b1001000001:out = 10'd192;
      10'b1001000010:out = 10'd192;
      10'b1001000011:out = 10'd193;
      10'b1001000100:out = 10'd193;
      10'b1001000101:out = 10'd193;
      10'b1001000110:out = 10'd194;
      10'b1001000111:out = 10'd194;
      10'b1001001000:out = 10'd194;
      10'b1001001001:out = 10'd195;
      10'b1001001010:out = 10'd195;
      10'b1001001011:out = 10'd195;
      10'b1001001100:out = 10'd196;
      10'b1001001101:out = 10'd196;
      10'b1001001110:out = 10'd196;
      10'b1001001111:out = 10'd197;
      10'b1001010000:out = 10'd197;
      10'b1001010001:out = 10'd197;
      10'b1001010010:out = 10'd198;
      10'b1001010011:out = 10'd198;
      10'b1001010100:out = 10'd198;
      10'b1001010101:out = 10'd199;
      10'b1001010110:out = 10'd199;
      10'b1001010111:out = 10'd199;
      10'b1001011000:out = 10'd200;
      10'b1001011001:out = 10'd200;
      10'b1001011010:out = 10'd200;
      10'b1001011011:out = 10'd201;
      10'b1001011100:out = 10'd201;
      10'b1001011101:out = 10'd201;
      10'b1001011110:out = 10'd202;
      10'b1001011111:out = 10'd202;
      10'b1001100000:out = 10'd202;
      10'b1001100001:out = 10'd203;
      10'b1001100010:out = 10'd203;
      10'b1001100011:out = 10'd203;
      10'b1001100100:out = 10'd204;
      10'b1001100101:out = 10'd204;
      10'b1001100110:out = 10'd204;
      10'b1001100111:out = 10'd205;
      10'b1001101000:out = 10'd205;
      10'b1001101001:out = 10'd205;
      10'b1001101010:out = 10'd206;
      10'b1001101011:out = 10'd206;
      10'b1001101100:out = 10'd206;
      10'b1001101101:out = 10'd207;
      10'b1001101110:out = 10'd207;
      10'b1001101111:out = 10'd207;
      10'b1001110000:out = 10'd208;
      10'b1001110001:out = 10'd208;
      10'b1001110010:out = 10'd208;
      10'b1001110011:out = 10'd209;
      10'b1001110100:out = 10'd209;
      10'b1001110101:out = 10'd209;
      10'b1001110110:out = 10'd210;
      10'b1001110111:out = 10'd210;
      10'b1001111000:out = 10'd210;
      10'b1001111001:out = 10'd211;
      10'b1001111010:out = 10'd211;
      10'b1001111011:out = 10'd211;
      10'b1001111100:out = 10'd212;
      10'b1001111101:out = 10'd212;
      10'b1001111110:out = 10'd212;
      10'b1001111111:out = 10'd213;
      10'b1010000000:out = 10'd213;
      10'b1010000001:out = 10'd213;
      10'b1010000010:out = 10'd214;
      10'b1010000011:out = 10'd214;
      10'b1010000100:out = 10'd214;
      10'b1010000101:out = 10'd215;
      10'b1010000110:out = 10'd215;
      10'b1010000111:out = 10'd215;
      10'b1010001000:out = 10'd216;
      10'b1010001001:out = 10'd216;
      10'b1010001010:out = 10'd216;
      10'b1010001011:out = 10'd217;
      10'b1010001100:out = 10'd217;
      10'b1010001101:out = 10'd217;
      10'b1010001110:out = 10'd218;
      10'b1010001111:out = 10'd218;
      10'b1010010000:out = 10'd218;
      10'b1010010001:out = 10'd219;
      10'b1010010010:out = 10'd219;
      10'b1010010011:out = 10'd219;
      10'b1010010100:out = 10'd220;
      10'b1010010101:out = 10'd220;
      10'b1010010110:out = 10'd220;
      10'b1010010111:out = 10'd221;
      10'b1010011000:out = 10'd221;
      10'b1010011001:out = 10'd221;
      10'b1010011010:out = 10'd222;
      10'b1010011011:out = 10'd222;
      10'b1010011100:out = 10'd222;
      10'b1010011101:out = 10'd223;
      10'b1010011110:out = 10'd223;
      10'b1010011111:out = 10'd223;
      10'b1010100000:out = 10'd224;
      10'b1010100001:out = 10'd224;
      10'b1010100010:out = 10'd224;
      10'b1010100011:out = 10'd225;
      10'b1010100100:out = 10'd225;
      10'b1010100101:out = 10'd225;
      10'b1010100110:out = 10'd226;
      10'b1010100111:out = 10'd226;
      10'b1010101000:out = 10'd226;
      10'b1010101001:out = 10'd227;
      10'b1010101010:out = 10'd227;
      10'b1010101011:out = 10'd227;
      10'b1010101100:out = 10'd228;
      10'b1010101101:out = 10'd228;
      10'b1010101110:out = 10'd228;
      10'b1010101111:out = 10'd229;
      10'b1010110000:out = 10'd229;
      10'b1010110001:out = 10'd229;
      10'b1010110010:out = 10'd230;
      10'b1010110011:out = 10'd230;
      10'b1010110100:out = 10'd230;
      10'b1010110101:out = 10'd231;
      10'b1010110110:out = 10'd231;
      10'b1010110111:out = 10'd231;
      10'b1010111000:out = 10'd232;
      10'b1010111001:out = 10'd232;
      10'b1010111010:out = 10'd232;
      10'b1010111011:out = 10'd233;
      10'b1010111100:out = 10'd233;
      10'b1010111101:out = 10'd233;
      10'b1010111110:out = 10'd234;
      10'b1010111111:out = 10'd234;
      10'b1011000000:out = 10'd234;
      10'b1011000001:out = 10'd235;
      10'b1011000010:out = 10'd235;
      10'b1011000011:out = 10'd235;
      10'b1011000100:out = 10'd236;
      10'b1011000101:out = 10'd236;
      10'b1011000110:out = 10'd236;
      10'b1011000111:out = 10'd237;
      10'b1011001000:out = 10'd237;
      10'b1011001001:out = 10'd237;
      10'b1011001010:out = 10'd238;
      10'b1011001011:out = 10'd238;
      10'b1011001100:out = 10'd238;
      10'b1011001101:out = 10'd239;
      10'b1011001110:out = 10'd239;
      10'b1011001111:out = 10'd239;
      10'b1011010000:out = 10'd240;
      10'b1011010001:out = 10'd240;
      10'b1011010010:out = 10'd240;
      10'b1011010011:out = 10'd241;
      10'b1011010100:out = 10'd241;
      10'b1011010101:out = 10'd241;
      10'b1011010110:out = 10'd242;
      10'b1011010111:out = 10'd242;
      10'b1011011000:out = 10'd242;
      10'b1011011001:out = 10'd243;
      10'b1011011010:out = 10'd243;
      10'b1011011011:out = 10'd243;
      10'b1011011100:out = 10'd244;
      10'b1011011101:out = 10'd244;
      10'b1011011110:out = 10'd244;
      10'b1011011111:out = 10'd245;
      10'b1011100000:out = 10'd245;
      10'b1011100001:out = 10'd245;
      10'b1011100010:out = 10'd246;
      10'b1011100011:out = 10'd246;
      10'b1011100100:out = 10'd246;
      10'b1011100101:out = 10'd247;
      10'b1011100110:out = 10'd247;
      10'b1011100111:out = 10'd247;
      10'b1011101000:out = 10'd248;
      10'b1011101001:out = 10'd248;
      10'b1011101010:out = 10'd248;
      10'b1011101011:out = 10'd249;
      10'b1011101100:out = 10'd249;
      10'b1011101101:out = 10'd249;
      10'b1011101110:out = 10'd250;
      10'b1011101111:out = 10'd250;
      10'b1011110000:out = 10'd250;
      10'b1011110001:out = 10'd251;
      10'b1011110010:out = 10'd251;
      10'b1011110011:out = 10'd251;
      10'b1011110100:out = 10'd252;
      10'b1011110101:out = 10'd252;
      10'b1011110110:out = 10'd252;
      10'b1011110111:out = 10'd253;
      10'b1011111000:out = 10'd253;
      10'b1011111001:out = 10'd253;
      10'b1011111010:out = 10'd254;
      10'b1011111011:out = 10'd254;
      10'b1011111100:out = 10'd254;
      10'b1011111101:out = 10'd255;
      10'b1011111110:out = 10'd255;
      10'b1011111111:out = 10'd255;
      10'b1100000000:out = 10'd256;
      10'b1100000001:out = 10'd256;
      10'b1100000010:out = 10'd256;
      10'b1100000011:out = 10'd257;
      10'b1100000100:out = 10'd257;
      10'b1100000101:out = 10'd257;
      10'b1100000110:out = 10'd258;
      10'b1100000111:out = 10'd258;
      10'b1100001000:out = 10'd258;
      10'b1100001001:out = 10'd259;
      10'b1100001010:out = 10'd259;
      10'b1100001011:out = 10'd259;
      10'b1100001100:out = 10'd260;
      10'b1100001101:out = 10'd260;
      10'b1100001110:out = 10'd260;
      10'b1100001111:out = 10'd261;
      10'b1100010000:out = 10'd261;
      10'b1100010001:out = 10'd261;
      10'b1100010010:out = 10'd262;
      10'b1100010011:out = 10'd262;
      10'b1100010100:out = 10'd262;
      10'b1100010101:out = 10'd263;
      10'b1100010110:out = 10'd263;
      10'b1100010111:out = 10'd263;
      10'b1100011000:out = 10'd264;
      10'b1100011001:out = 10'd264;
      10'b1100011010:out = 10'd264;
      10'b1100011011:out = 10'd265;
      10'b1100011100:out = 10'd265;
      10'b1100011101:out = 10'd265;
      10'b1100011110:out = 10'd266;
      10'b1100011111:out = 10'd266;
      10'b1100100000:out = 10'd266;
      10'b1100100001:out = 10'd267;
      10'b1100100010:out = 10'd267;
      10'b1100100011:out = 10'd267;
      10'b1100100100:out = 10'd268;
      10'b1100100101:out = 10'd268;
      10'b1100100110:out = 10'd268;
      10'b1100100111:out = 10'd269;
      10'b1100101000:out = 10'd269;
      10'b1100101001:out = 10'd269;
      10'b1100101010:out = 10'd270;
      10'b1100101011:out = 10'd270;
      10'b1100101100:out = 10'd270;
      10'b1100101101:out = 10'd271;
      10'b1100101110:out = 10'd271;
      10'b1100101111:out = 10'd271;
      10'b1100110000:out = 10'd272;
      10'b1100110001:out = 10'd272;
      10'b1100110010:out = 10'd272;
      10'b1100110011:out = 10'd273;
      10'b1100110100:out = 10'd273;
      10'b1100110101:out = 10'd273;
      10'b1100110110:out = 10'd274;
      10'b1100110111:out = 10'd274;
      10'b1100111000:out = 10'd274;
      10'b1100111001:out = 10'd275;
      10'b1100111010:out = 10'd275;
      10'b1100111011:out = 10'd275;
      10'b1100111100:out = 10'd276;
      10'b1100111101:out = 10'd276;
      10'b1100111110:out = 10'd276;
      10'b1100111111:out = 10'd277;
      10'b1101000000:out = 10'd277;
      10'b1101000001:out = 10'd277;
      10'b1101000010:out = 10'd278;
      10'b1101000011:out = 10'd278;
      10'b1101000100:out = 10'd278;
      10'b1101000101:out = 10'd279;
      10'b1101000110:out = 10'd279;
      10'b1101000111:out = 10'd279;
      10'b1101001000:out = 10'd280;
      10'b1101001001:out = 10'd280;
      10'b1101001010:out = 10'd280;
      10'b1101001011:out = 10'd281;
      10'b1101001100:out = 10'd281;
      10'b1101001101:out = 10'd281;
      10'b1101001110:out = 10'd282;
      10'b1101001111:out = 10'd282;
      10'b1101010000:out = 10'd282;
      10'b1101010001:out = 10'd283;
      10'b1101010010:out = 10'd283;
      10'b1101010011:out = 10'd283;
      10'b1101010100:out = 10'd284;
      10'b1101010101:out = 10'd284;
      10'b1101010110:out = 10'd284;
      10'b1101010111:out = 10'd285;
      10'b1101011000:out = 10'd285;
      10'b1101011001:out = 10'd285;
      10'b1101011010:out = 10'd286;
      10'b1101011011:out = 10'd286;
      10'b1101011100:out = 10'd286;
      10'b1101011101:out = 10'd287;
      10'b1101011110:out = 10'd287;
      10'b1101011111:out = 10'd287;
      10'b1101100000:out = 10'd288;
      10'b1101100001:out = 10'd288;
      10'b1101100010:out = 10'd288;
      10'b1101100011:out = 10'd289;
      10'b1101100100:out = 10'd289;
      10'b1101100101:out = 10'd289;
      10'b1101100110:out = 10'd290;
      10'b1101100111:out = 10'd290;
      10'b1101101000:out = 10'd290;
      10'b1101101001:out = 10'd291;
      10'b1101101010:out = 10'd291;
      10'b1101101011:out = 10'd291;
      10'b1101101100:out = 10'd292;
      10'b1101101101:out = 10'd292;
      10'b1101101110:out = 10'd292;
      10'b1101101111:out = 10'd293;
      10'b1101110000:out = 10'd293;
      10'b1101110001:out = 10'd293;
      10'b1101110010:out = 10'd294;
      10'b1101110011:out = 10'd294;
      10'b1101110100:out = 10'd294;
      10'b1101110101:out = 10'd295;
      10'b1101110110:out = 10'd295;
      10'b1101110111:out = 10'd295;
      10'b1101111000:out = 10'd296;
      10'b1101111001:out = 10'd296;
      10'b1101111010:out = 10'd296;
      10'b1101111011:out = 10'd297;
      10'b1101111100:out = 10'd297;
      10'b1101111101:out = 10'd297;
      10'b1101111110:out = 10'd298;
      10'b1101111111:out = 10'd298;
      10'b1110000000:out = 10'd298;
      10'b1110000001:out = 10'd299;
      10'b1110000010:out = 10'd299;
      10'b1110000011:out = 10'd299;
      10'b1110000100:out = 10'd300;
      10'b1110000101:out = 10'd300;
      10'b1110000110:out = 10'd300;
      10'b1110000111:out = 10'd301;
      10'b1110001000:out = 10'd301;
      10'b1110001001:out = 10'd301;
      10'b1110001010:out = 10'd302;
      10'b1110001011:out = 10'd302;
      10'b1110001100:out = 10'd302;
      10'b1110001101:out = 10'd303;
      10'b1110001110:out = 10'd303;
      10'b1110001111:out = 10'd303;
      10'b1110010000:out = 10'd304;
      10'b1110010001:out = 10'd304;
      10'b1110010010:out = 10'd304;
      10'b1110010011:out = 10'd305;
      10'b1110010100:out = 10'd305;
      10'b1110010101:out = 10'd305;
      10'b1110010110:out = 10'd306;
      10'b1110010111:out = 10'd306;
      10'b1110011000:out = 10'd306;
      10'b1110011001:out = 10'd307;
      10'b1110011010:out = 10'd307;
      10'b1110011011:out = 10'd307;
      10'b1110011100:out = 10'd308;
      10'b1110011101:out = 10'd308;
      10'b1110011110:out = 10'd308;
      10'b1110011111:out = 10'd309;
      10'b1110100000:out = 10'd309;
      10'b1110100001:out = 10'd309;
      10'b1110100010:out = 10'd310;
      10'b1110100011:out = 10'd310;
      10'b1110100100:out = 10'd310;
      10'b1110100101:out = 10'd311;
      10'b1110100110:out = 10'd311;
      10'b1110100111:out = 10'd311;
      10'b1110101000:out = 10'd312;
      10'b1110101001:out = 10'd312;
      10'b1110101010:out = 10'd312;
      10'b1110101011:out = 10'd313;
      10'b1110101100:out = 10'd313;
      10'b1110101101:out = 10'd313;
      10'b1110101110:out = 10'd314;
      10'b1110101111:out = 10'd314;
      10'b1110110000:out = 10'd314;
      10'b1110110001:out = 10'd315;
      10'b1110110010:out = 10'd315;
      10'b1110110011:out = 10'd315;
      10'b1110110100:out = 10'd316;
      10'b1110110101:out = 10'd316;
      10'b1110110110:out = 10'd316;
      10'b1110110111:out = 10'd317;
      10'b1110111000:out = 10'd317;
      10'b1110111001:out = 10'd317;
      10'b1110111010:out = 10'd318;
      10'b1110111011:out = 10'd318;
      10'b1110111100:out = 10'd318;
      10'b1110111101:out = 10'd319;
      10'b1110111110:out = 10'd319;
      10'b1110111111:out = 10'd319;
      10'b1111000000:out = 10'd320;
      10'b1111000001:out = 10'd320;
      10'b1111000010:out = 10'd320;
      10'b1111000011:out = 10'd321;
      10'b1111000100:out = 10'd321;
      10'b1111000101:out = 10'd321;
      10'b1111000110:out = 10'd322;
      10'b1111000111:out = 10'd322;
      10'b1111001000:out = 10'd322;
      10'b1111001001:out = 10'd323;
      10'b1111001010:out = 10'd323;
      10'b1111001011:out = 10'd323;
      10'b1111001100:out = 10'd324;
      10'b1111001101:out = 10'd324;
      10'b1111001110:out = 10'd324;
      10'b1111001111:out = 10'd325;
      10'b1111010000:out = 10'd325;
      10'b1111010001:out = 10'd325;
      10'b1111010010:out = 10'd326;
      10'b1111010011:out = 10'd326;
      10'b1111010100:out = 10'd326;
      10'b1111010101:out = 10'd327;
      10'b1111010110:out = 10'd327;
      10'b1111010111:out = 10'd327;
      10'b1111011000:out = 10'd328;
      10'b1111011001:out = 10'd328;
      10'b1111011010:out = 10'd328;
      10'b1111011011:out = 10'd329;
      10'b1111011100:out = 10'd329;
      10'b1111011101:out = 10'd329;
      10'b1111011110:out = 10'd330;
      10'b1111011111:out = 10'd330;
      10'b1111100000:out = 10'd330;
      10'b1111100001:out = 10'd331;
      10'b1111100010:out = 10'd331;
      10'b1111100011:out = 10'd331;
      10'b1111100100:out = 10'd332;
      10'b1111100101:out = 10'd332;
      10'b1111100110:out = 10'd332;
      10'b1111100111:out = 10'd333;
      10'b1111101000:out = 10'd333;
      10'b1111101001:out = 10'd333;
      10'b1111101010:out = 10'd334;
      10'b1111101011:out = 10'd334;
      10'b1111101100:out = 10'd334;
      10'b1111101101:out = 10'd335;
      10'b1111101110:out = 10'd335;
      10'b1111101111:out = 10'd335;
      10'b1111110000:out = 10'd336;
      10'b1111110001:out = 10'd336;
      10'b1111110010:out = 10'd336;
      10'b1111110011:out = 10'd337;
      10'b1111110100:out = 10'd337;
      10'b1111110101:out = 10'd337;
      10'b1111110110:out = 10'd338;
      10'b1111110111:out = 10'd338;
      10'b1111111000:out = 10'd338;
      10'b1111111001:out = 10'd339;
      10'b1111111010:out = 10'd339;
      10'b1111111011:out = 10'd339;
      10'b1111111100:out = 10'd340;
      10'b1111111101:out = 10'd340;
      10'b1111111110:out = 10'd340;
      10'b1111111111:out = 10'd341;
    endcase
  end
endmodule

