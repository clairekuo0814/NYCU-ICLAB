# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : MEM5x5
#       Words            : 416
#       Bits             : 8
#       Byte-Write       : 1
#       Aspect Ratio     : 2
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2023/11/28 01:36:31
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO MEM5x5
CLASS BLOCK ;
FOREIGN MEM5x5 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 316.200 BY 201.040 ;
SYMMETRY x y r90 ;
SITE core_5040 ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 315.080 188.500 316.200 191.740 ;
  LAYER metal3 ;
  RECT 315.080 188.500 316.200 191.740 ;
  LAYER metal2 ;
  RECT 315.080 188.500 316.200 191.740 ;
  LAYER metal1 ;
  RECT 315.080 188.500 316.200 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 180.660 316.200 183.900 ;
  LAYER metal3 ;
  RECT 315.080 180.660 316.200 183.900 ;
  LAYER metal2 ;
  RECT 315.080 180.660 316.200 183.900 ;
  LAYER metal1 ;
  RECT 315.080 180.660 316.200 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 172.820 316.200 176.060 ;
  LAYER metal3 ;
  RECT 315.080 172.820 316.200 176.060 ;
  LAYER metal2 ;
  RECT 315.080 172.820 316.200 176.060 ;
  LAYER metal1 ;
  RECT 315.080 172.820 316.200 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 164.980 316.200 168.220 ;
  LAYER metal3 ;
  RECT 315.080 164.980 316.200 168.220 ;
  LAYER metal2 ;
  RECT 315.080 164.980 316.200 168.220 ;
  LAYER metal1 ;
  RECT 315.080 164.980 316.200 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 125.780 316.200 129.020 ;
  LAYER metal3 ;
  RECT 315.080 125.780 316.200 129.020 ;
  LAYER metal2 ;
  RECT 315.080 125.780 316.200 129.020 ;
  LAYER metal1 ;
  RECT 315.080 125.780 316.200 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 117.940 316.200 121.180 ;
  LAYER metal3 ;
  RECT 315.080 117.940 316.200 121.180 ;
  LAYER metal2 ;
  RECT 315.080 117.940 316.200 121.180 ;
  LAYER metal1 ;
  RECT 315.080 117.940 316.200 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 110.100 316.200 113.340 ;
  LAYER metal3 ;
  RECT 315.080 110.100 316.200 113.340 ;
  LAYER metal2 ;
  RECT 315.080 110.100 316.200 113.340 ;
  LAYER metal1 ;
  RECT 315.080 110.100 316.200 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 102.260 316.200 105.500 ;
  LAYER metal3 ;
  RECT 315.080 102.260 316.200 105.500 ;
  LAYER metal2 ;
  RECT 315.080 102.260 316.200 105.500 ;
  LAYER metal1 ;
  RECT 315.080 102.260 316.200 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 94.420 316.200 97.660 ;
  LAYER metal3 ;
  RECT 315.080 94.420 316.200 97.660 ;
  LAYER metal2 ;
  RECT 315.080 94.420 316.200 97.660 ;
  LAYER metal1 ;
  RECT 315.080 94.420 316.200 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 86.580 316.200 89.820 ;
  LAYER metal3 ;
  RECT 315.080 86.580 316.200 89.820 ;
  LAYER metal2 ;
  RECT 315.080 86.580 316.200 89.820 ;
  LAYER metal1 ;
  RECT 315.080 86.580 316.200 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 47.380 316.200 50.620 ;
  LAYER metal3 ;
  RECT 315.080 47.380 316.200 50.620 ;
  LAYER metal2 ;
  RECT 315.080 47.380 316.200 50.620 ;
  LAYER metal1 ;
  RECT 315.080 47.380 316.200 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 39.540 316.200 42.780 ;
  LAYER metal3 ;
  RECT 315.080 39.540 316.200 42.780 ;
  LAYER metal2 ;
  RECT 315.080 39.540 316.200 42.780 ;
  LAYER metal1 ;
  RECT 315.080 39.540 316.200 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 31.700 316.200 34.940 ;
  LAYER metal3 ;
  RECT 315.080 31.700 316.200 34.940 ;
  LAYER metal2 ;
  RECT 315.080 31.700 316.200 34.940 ;
  LAYER metal1 ;
  RECT 315.080 31.700 316.200 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 23.860 316.200 27.100 ;
  LAYER metal3 ;
  RECT 315.080 23.860 316.200 27.100 ;
  LAYER metal2 ;
  RECT 315.080 23.860 316.200 27.100 ;
  LAYER metal1 ;
  RECT 315.080 23.860 316.200 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 16.020 316.200 19.260 ;
  LAYER metal3 ;
  RECT 315.080 16.020 316.200 19.260 ;
  LAYER metal2 ;
  RECT 315.080 16.020 316.200 19.260 ;
  LAYER metal1 ;
  RECT 315.080 16.020 316.200 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 8.180 316.200 11.420 ;
  LAYER metal3 ;
  RECT 315.080 8.180 316.200 11.420 ;
  LAYER metal2 ;
  RECT 315.080 8.180 316.200 11.420 ;
  LAYER metal1 ;
  RECT 315.080 8.180 316.200 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 302.960 199.920 306.500 201.040 ;
  LAYER metal3 ;
  RECT 302.960 199.920 306.500 201.040 ;
  LAYER metal2 ;
  RECT 302.960 199.920 306.500 201.040 ;
  LAYER metal1 ;
  RECT 302.960 199.920 306.500 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 294.280 199.920 297.820 201.040 ;
  LAYER metal3 ;
  RECT 294.280 199.920 297.820 201.040 ;
  LAYER metal2 ;
  RECT 294.280 199.920 297.820 201.040 ;
  LAYER metal1 ;
  RECT 294.280 199.920 297.820 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 285.600 199.920 289.140 201.040 ;
  LAYER metal3 ;
  RECT 285.600 199.920 289.140 201.040 ;
  LAYER metal2 ;
  RECT 285.600 199.920 289.140 201.040 ;
  LAYER metal1 ;
  RECT 285.600 199.920 289.140 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 276.920 199.920 280.460 201.040 ;
  LAYER metal3 ;
  RECT 276.920 199.920 280.460 201.040 ;
  LAYER metal2 ;
  RECT 276.920 199.920 280.460 201.040 ;
  LAYER metal1 ;
  RECT 276.920 199.920 280.460 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 268.240 199.920 271.780 201.040 ;
  LAYER metal3 ;
  RECT 268.240 199.920 271.780 201.040 ;
  LAYER metal2 ;
  RECT 268.240 199.920 271.780 201.040 ;
  LAYER metal1 ;
  RECT 268.240 199.920 271.780 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 224.840 199.920 228.380 201.040 ;
  LAYER metal3 ;
  RECT 224.840 199.920 228.380 201.040 ;
  LAYER metal2 ;
  RECT 224.840 199.920 228.380 201.040 ;
  LAYER metal1 ;
  RECT 224.840 199.920 228.380 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 216.160 199.920 219.700 201.040 ;
  LAYER metal3 ;
  RECT 216.160 199.920 219.700 201.040 ;
  LAYER metal2 ;
  RECT 216.160 199.920 219.700 201.040 ;
  LAYER metal1 ;
  RECT 216.160 199.920 219.700 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 207.480 199.920 211.020 201.040 ;
  LAYER metal3 ;
  RECT 207.480 199.920 211.020 201.040 ;
  LAYER metal2 ;
  RECT 207.480 199.920 211.020 201.040 ;
  LAYER metal1 ;
  RECT 207.480 199.920 211.020 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.800 199.920 202.340 201.040 ;
  LAYER metal3 ;
  RECT 198.800 199.920 202.340 201.040 ;
  LAYER metal2 ;
  RECT 198.800 199.920 202.340 201.040 ;
  LAYER metal1 ;
  RECT 198.800 199.920 202.340 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.120 199.920 193.660 201.040 ;
  LAYER metal3 ;
  RECT 190.120 199.920 193.660 201.040 ;
  LAYER metal2 ;
  RECT 190.120 199.920 193.660 201.040 ;
  LAYER metal1 ;
  RECT 190.120 199.920 193.660 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 181.440 199.920 184.980 201.040 ;
  LAYER metal3 ;
  RECT 181.440 199.920 184.980 201.040 ;
  LAYER metal2 ;
  RECT 181.440 199.920 184.980 201.040 ;
  LAYER metal1 ;
  RECT 181.440 199.920 184.980 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 138.040 199.920 141.580 201.040 ;
  LAYER metal3 ;
  RECT 138.040 199.920 141.580 201.040 ;
  LAYER metal2 ;
  RECT 138.040 199.920 141.580 201.040 ;
  LAYER metal1 ;
  RECT 138.040 199.920 141.580 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 129.360 199.920 132.900 201.040 ;
  LAYER metal3 ;
  RECT 129.360 199.920 132.900 201.040 ;
  LAYER metal2 ;
  RECT 129.360 199.920 132.900 201.040 ;
  LAYER metal1 ;
  RECT 129.360 199.920 132.900 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 120.680 199.920 124.220 201.040 ;
  LAYER metal3 ;
  RECT 120.680 199.920 124.220 201.040 ;
  LAYER metal2 ;
  RECT 120.680 199.920 124.220 201.040 ;
  LAYER metal1 ;
  RECT 120.680 199.920 124.220 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 112.000 199.920 115.540 201.040 ;
  LAYER metal3 ;
  RECT 112.000 199.920 115.540 201.040 ;
  LAYER metal2 ;
  RECT 112.000 199.920 115.540 201.040 ;
  LAYER metal1 ;
  RECT 112.000 199.920 115.540 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 103.320 199.920 106.860 201.040 ;
  LAYER metal3 ;
  RECT 103.320 199.920 106.860 201.040 ;
  LAYER metal2 ;
  RECT 103.320 199.920 106.860 201.040 ;
  LAYER metal1 ;
  RECT 103.320 199.920 106.860 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 94.640 199.920 98.180 201.040 ;
  LAYER metal3 ;
  RECT 94.640 199.920 98.180 201.040 ;
  LAYER metal2 ;
  RECT 94.640 199.920 98.180 201.040 ;
  LAYER metal1 ;
  RECT 94.640 199.920 98.180 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 51.240 199.920 54.780 201.040 ;
  LAYER metal3 ;
  RECT 51.240 199.920 54.780 201.040 ;
  LAYER metal2 ;
  RECT 51.240 199.920 54.780 201.040 ;
  LAYER metal1 ;
  RECT 51.240 199.920 54.780 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 42.560 199.920 46.100 201.040 ;
  LAYER metal3 ;
  RECT 42.560 199.920 46.100 201.040 ;
  LAYER metal2 ;
  RECT 42.560 199.920 46.100 201.040 ;
  LAYER metal1 ;
  RECT 42.560 199.920 46.100 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.880 199.920 37.420 201.040 ;
  LAYER metal3 ;
  RECT 33.880 199.920 37.420 201.040 ;
  LAYER metal2 ;
  RECT 33.880 199.920 37.420 201.040 ;
  LAYER metal1 ;
  RECT 33.880 199.920 37.420 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.200 199.920 28.740 201.040 ;
  LAYER metal3 ;
  RECT 25.200 199.920 28.740 201.040 ;
  LAYER metal2 ;
  RECT 25.200 199.920 28.740 201.040 ;
  LAYER metal1 ;
  RECT 25.200 199.920 28.740 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 16.520 199.920 20.060 201.040 ;
  LAYER metal3 ;
  RECT 16.520 199.920 20.060 201.040 ;
  LAYER metal2 ;
  RECT 16.520 199.920 20.060 201.040 ;
  LAYER metal1 ;
  RECT 16.520 199.920 20.060 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.840 199.920 11.380 201.040 ;
  LAYER metal3 ;
  RECT 7.840 199.920 11.380 201.040 ;
  LAYER metal2 ;
  RECT 7.840 199.920 11.380 201.040 ;
  LAYER metal1 ;
  RECT 7.840 199.920 11.380 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 301.100 0.000 304.640 1.120 ;
  LAYER metal3 ;
  RECT 301.100 0.000 304.640 1.120 ;
  LAYER metal2 ;
  RECT 301.100 0.000 304.640 1.120 ;
  LAYER metal1 ;
  RECT 301.100 0.000 304.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 292.420 0.000 295.960 1.120 ;
  LAYER metal3 ;
  RECT 292.420 0.000 295.960 1.120 ;
  LAYER metal2 ;
  RECT 292.420 0.000 295.960 1.120 ;
  LAYER metal1 ;
  RECT 292.420 0.000 295.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 231.660 0.000 235.200 1.120 ;
  LAYER metal3 ;
  RECT 231.660 0.000 235.200 1.120 ;
  LAYER metal2 ;
  RECT 231.660 0.000 235.200 1.120 ;
  LAYER metal1 ;
  RECT 231.660 0.000 235.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 222.980 0.000 226.520 1.120 ;
  LAYER metal3 ;
  RECT 222.980 0.000 226.520 1.120 ;
  LAYER metal2 ;
  RECT 222.980 0.000 226.520 1.120 ;
  LAYER metal1 ;
  RECT 222.980 0.000 226.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 209.960 0.000 213.500 1.120 ;
  LAYER metal3 ;
  RECT 209.960 0.000 213.500 1.120 ;
  LAYER metal2 ;
  RECT 209.960 0.000 213.500 1.120 ;
  LAYER metal1 ;
  RECT 209.960 0.000 213.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 174.000 0.000 177.540 1.120 ;
  LAYER metal3 ;
  RECT 174.000 0.000 177.540 1.120 ;
  LAYER metal2 ;
  RECT 174.000 0.000 177.540 1.120 ;
  LAYER metal1 ;
  RECT 174.000 0.000 177.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 165.320 0.000 168.860 1.120 ;
  LAYER metal3 ;
  RECT 165.320 0.000 168.860 1.120 ;
  LAYER metal2 ;
  RECT 165.320 0.000 168.860 1.120 ;
  LAYER metal1 ;
  RECT 165.320 0.000 168.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 143.620 0.000 147.160 1.120 ;
  LAYER metal3 ;
  RECT 143.620 0.000 147.160 1.120 ;
  LAYER metal2 ;
  RECT 143.620 0.000 147.160 1.120 ;
  LAYER metal1 ;
  RECT 143.620 0.000 147.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal3 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal2 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal1 ;
  RECT 61.780 0.000 65.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal3 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal2 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal1 ;
  RECT 53.100 0.000 56.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal3 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal2 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal1 ;
  RECT 44.420 0.000 47.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 315.080 184.580 316.200 187.820 ;
  LAYER metal3 ;
  RECT 315.080 184.580 316.200 187.820 ;
  LAYER metal2 ;
  RECT 315.080 184.580 316.200 187.820 ;
  LAYER metal1 ;
  RECT 315.080 184.580 316.200 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 176.740 316.200 179.980 ;
  LAYER metal3 ;
  RECT 315.080 176.740 316.200 179.980 ;
  LAYER metal2 ;
  RECT 315.080 176.740 316.200 179.980 ;
  LAYER metal1 ;
  RECT 315.080 176.740 316.200 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 168.900 316.200 172.140 ;
  LAYER metal3 ;
  RECT 315.080 168.900 316.200 172.140 ;
  LAYER metal2 ;
  RECT 315.080 168.900 316.200 172.140 ;
  LAYER metal1 ;
  RECT 315.080 168.900 316.200 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 129.700 316.200 132.940 ;
  LAYER metal3 ;
  RECT 315.080 129.700 316.200 132.940 ;
  LAYER metal2 ;
  RECT 315.080 129.700 316.200 132.940 ;
  LAYER metal1 ;
  RECT 315.080 129.700 316.200 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 121.860 316.200 125.100 ;
  LAYER metal3 ;
  RECT 315.080 121.860 316.200 125.100 ;
  LAYER metal2 ;
  RECT 315.080 121.860 316.200 125.100 ;
  LAYER metal1 ;
  RECT 315.080 121.860 316.200 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 114.020 316.200 117.260 ;
  LAYER metal3 ;
  RECT 315.080 114.020 316.200 117.260 ;
  LAYER metal2 ;
  RECT 315.080 114.020 316.200 117.260 ;
  LAYER metal1 ;
  RECT 315.080 114.020 316.200 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 106.180 316.200 109.420 ;
  LAYER metal3 ;
  RECT 315.080 106.180 316.200 109.420 ;
  LAYER metal2 ;
  RECT 315.080 106.180 316.200 109.420 ;
  LAYER metal1 ;
  RECT 315.080 106.180 316.200 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 98.340 316.200 101.580 ;
  LAYER metal3 ;
  RECT 315.080 98.340 316.200 101.580 ;
  LAYER metal2 ;
  RECT 315.080 98.340 316.200 101.580 ;
  LAYER metal1 ;
  RECT 315.080 98.340 316.200 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 90.500 316.200 93.740 ;
  LAYER metal3 ;
  RECT 315.080 90.500 316.200 93.740 ;
  LAYER metal2 ;
  RECT 315.080 90.500 316.200 93.740 ;
  LAYER metal1 ;
  RECT 315.080 90.500 316.200 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 51.300 316.200 54.540 ;
  LAYER metal3 ;
  RECT 315.080 51.300 316.200 54.540 ;
  LAYER metal2 ;
  RECT 315.080 51.300 316.200 54.540 ;
  LAYER metal1 ;
  RECT 315.080 51.300 316.200 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 43.460 316.200 46.700 ;
  LAYER metal3 ;
  RECT 315.080 43.460 316.200 46.700 ;
  LAYER metal2 ;
  RECT 315.080 43.460 316.200 46.700 ;
  LAYER metal1 ;
  RECT 315.080 43.460 316.200 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 35.620 316.200 38.860 ;
  LAYER metal3 ;
  RECT 315.080 35.620 316.200 38.860 ;
  LAYER metal2 ;
  RECT 315.080 35.620 316.200 38.860 ;
  LAYER metal1 ;
  RECT 315.080 35.620 316.200 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 27.780 316.200 31.020 ;
  LAYER metal3 ;
  RECT 315.080 27.780 316.200 31.020 ;
  LAYER metal2 ;
  RECT 315.080 27.780 316.200 31.020 ;
  LAYER metal1 ;
  RECT 315.080 27.780 316.200 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 19.940 316.200 23.180 ;
  LAYER metal3 ;
  RECT 315.080 19.940 316.200 23.180 ;
  LAYER metal2 ;
  RECT 315.080 19.940 316.200 23.180 ;
  LAYER metal1 ;
  RECT 315.080 19.940 316.200 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.080 12.100 316.200 15.340 ;
  LAYER metal3 ;
  RECT 315.080 12.100 316.200 15.340 ;
  LAYER metal2 ;
  RECT 315.080 12.100 316.200 15.340 ;
  LAYER metal1 ;
  RECT 315.080 12.100 316.200 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 298.620 199.920 302.160 201.040 ;
  LAYER metal3 ;
  RECT 298.620 199.920 302.160 201.040 ;
  LAYER metal2 ;
  RECT 298.620 199.920 302.160 201.040 ;
  LAYER metal1 ;
  RECT 298.620 199.920 302.160 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 289.940 199.920 293.480 201.040 ;
  LAYER metal3 ;
  RECT 289.940 199.920 293.480 201.040 ;
  LAYER metal2 ;
  RECT 289.940 199.920 293.480 201.040 ;
  LAYER metal1 ;
  RECT 289.940 199.920 293.480 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 281.260 199.920 284.800 201.040 ;
  LAYER metal3 ;
  RECT 281.260 199.920 284.800 201.040 ;
  LAYER metal2 ;
  RECT 281.260 199.920 284.800 201.040 ;
  LAYER metal1 ;
  RECT 281.260 199.920 284.800 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 272.580 199.920 276.120 201.040 ;
  LAYER metal3 ;
  RECT 272.580 199.920 276.120 201.040 ;
  LAYER metal2 ;
  RECT 272.580 199.920 276.120 201.040 ;
  LAYER metal1 ;
  RECT 272.580 199.920 276.120 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.180 199.920 232.720 201.040 ;
  LAYER metal3 ;
  RECT 229.180 199.920 232.720 201.040 ;
  LAYER metal2 ;
  RECT 229.180 199.920 232.720 201.040 ;
  LAYER metal1 ;
  RECT 229.180 199.920 232.720 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 220.500 199.920 224.040 201.040 ;
  LAYER metal3 ;
  RECT 220.500 199.920 224.040 201.040 ;
  LAYER metal2 ;
  RECT 220.500 199.920 224.040 201.040 ;
  LAYER metal1 ;
  RECT 220.500 199.920 224.040 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 211.820 199.920 215.360 201.040 ;
  LAYER metal3 ;
  RECT 211.820 199.920 215.360 201.040 ;
  LAYER metal2 ;
  RECT 211.820 199.920 215.360 201.040 ;
  LAYER metal1 ;
  RECT 211.820 199.920 215.360 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 203.140 199.920 206.680 201.040 ;
  LAYER metal3 ;
  RECT 203.140 199.920 206.680 201.040 ;
  LAYER metal2 ;
  RECT 203.140 199.920 206.680 201.040 ;
  LAYER metal1 ;
  RECT 203.140 199.920 206.680 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 194.460 199.920 198.000 201.040 ;
  LAYER metal3 ;
  RECT 194.460 199.920 198.000 201.040 ;
  LAYER metal2 ;
  RECT 194.460 199.920 198.000 201.040 ;
  LAYER metal1 ;
  RECT 194.460 199.920 198.000 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 185.780 199.920 189.320 201.040 ;
  LAYER metal3 ;
  RECT 185.780 199.920 189.320 201.040 ;
  LAYER metal2 ;
  RECT 185.780 199.920 189.320 201.040 ;
  LAYER metal1 ;
  RECT 185.780 199.920 189.320 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.380 199.920 145.920 201.040 ;
  LAYER metal3 ;
  RECT 142.380 199.920 145.920 201.040 ;
  LAYER metal2 ;
  RECT 142.380 199.920 145.920 201.040 ;
  LAYER metal1 ;
  RECT 142.380 199.920 145.920 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 133.700 199.920 137.240 201.040 ;
  LAYER metal3 ;
  RECT 133.700 199.920 137.240 201.040 ;
  LAYER metal2 ;
  RECT 133.700 199.920 137.240 201.040 ;
  LAYER metal1 ;
  RECT 133.700 199.920 137.240 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.020 199.920 128.560 201.040 ;
  LAYER metal3 ;
  RECT 125.020 199.920 128.560 201.040 ;
  LAYER metal2 ;
  RECT 125.020 199.920 128.560 201.040 ;
  LAYER metal1 ;
  RECT 125.020 199.920 128.560 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 116.340 199.920 119.880 201.040 ;
  LAYER metal3 ;
  RECT 116.340 199.920 119.880 201.040 ;
  LAYER metal2 ;
  RECT 116.340 199.920 119.880 201.040 ;
  LAYER metal1 ;
  RECT 116.340 199.920 119.880 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.660 199.920 111.200 201.040 ;
  LAYER metal3 ;
  RECT 107.660 199.920 111.200 201.040 ;
  LAYER metal2 ;
  RECT 107.660 199.920 111.200 201.040 ;
  LAYER metal1 ;
  RECT 107.660 199.920 111.200 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 98.980 199.920 102.520 201.040 ;
  LAYER metal3 ;
  RECT 98.980 199.920 102.520 201.040 ;
  LAYER metal2 ;
  RECT 98.980 199.920 102.520 201.040 ;
  LAYER metal1 ;
  RECT 98.980 199.920 102.520 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 55.580 199.920 59.120 201.040 ;
  LAYER metal3 ;
  RECT 55.580 199.920 59.120 201.040 ;
  LAYER metal2 ;
  RECT 55.580 199.920 59.120 201.040 ;
  LAYER metal1 ;
  RECT 55.580 199.920 59.120 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 46.900 199.920 50.440 201.040 ;
  LAYER metal3 ;
  RECT 46.900 199.920 50.440 201.040 ;
  LAYER metal2 ;
  RECT 46.900 199.920 50.440 201.040 ;
  LAYER metal1 ;
  RECT 46.900 199.920 50.440 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 38.220 199.920 41.760 201.040 ;
  LAYER metal3 ;
  RECT 38.220 199.920 41.760 201.040 ;
  LAYER metal2 ;
  RECT 38.220 199.920 41.760 201.040 ;
  LAYER metal1 ;
  RECT 38.220 199.920 41.760 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.540 199.920 33.080 201.040 ;
  LAYER metal3 ;
  RECT 29.540 199.920 33.080 201.040 ;
  LAYER metal2 ;
  RECT 29.540 199.920 33.080 201.040 ;
  LAYER metal1 ;
  RECT 29.540 199.920 33.080 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 20.860 199.920 24.400 201.040 ;
  LAYER metal3 ;
  RECT 20.860 199.920 24.400 201.040 ;
  LAYER metal2 ;
  RECT 20.860 199.920 24.400 201.040 ;
  LAYER metal1 ;
  RECT 20.860 199.920 24.400 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.180 199.920 15.720 201.040 ;
  LAYER metal3 ;
  RECT 12.180 199.920 15.720 201.040 ;
  LAYER metal2 ;
  RECT 12.180 199.920 15.720 201.040 ;
  LAYER metal1 ;
  RECT 12.180 199.920 15.720 201.040 ;
 END
 PORT
  LAYER metal4 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal3 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal2 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal1 ;
  RECT 296.760 0.000 300.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 236.000 0.000 239.540 1.120 ;
  LAYER metal3 ;
  RECT 236.000 0.000 239.540 1.120 ;
  LAYER metal2 ;
  RECT 236.000 0.000 239.540 1.120 ;
  LAYER metal1 ;
  RECT 236.000 0.000 239.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 227.320 0.000 230.860 1.120 ;
  LAYER metal3 ;
  RECT 227.320 0.000 230.860 1.120 ;
  LAYER metal2 ;
  RECT 227.320 0.000 230.860 1.120 ;
  LAYER metal1 ;
  RECT 227.320 0.000 230.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 218.640 0.000 222.180 1.120 ;
  LAYER metal3 ;
  RECT 218.640 0.000 222.180 1.120 ;
  LAYER metal2 ;
  RECT 218.640 0.000 222.180 1.120 ;
  LAYER metal1 ;
  RECT 218.640 0.000 222.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 196.940 0.000 200.480 1.120 ;
  LAYER metal3 ;
  RECT 196.940 0.000 200.480 1.120 ;
  LAYER metal2 ;
  RECT 196.940 0.000 200.480 1.120 ;
  LAYER metal1 ;
  RECT 196.940 0.000 200.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 169.660 0.000 173.200 1.120 ;
  LAYER metal3 ;
  RECT 169.660 0.000 173.200 1.120 ;
  LAYER metal2 ;
  RECT 169.660 0.000 173.200 1.120 ;
  LAYER metal1 ;
  RECT 169.660 0.000 173.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 160.980 0.000 164.520 1.120 ;
  LAYER metal3 ;
  RECT 160.980 0.000 164.520 1.120 ;
  LAYER metal2 ;
  RECT 160.980 0.000 164.520 1.120 ;
  LAYER metal1 ;
  RECT 160.980 0.000 164.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal3 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal2 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal1 ;
  RECT 57.440 0.000 60.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal3 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal2 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal1 ;
  RECT 48.760 0.000 52.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal3 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal2 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal1 ;
  RECT 40.080 0.000 43.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER metal4 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER metal3 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER metal2 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER metal1 ;
  RECT 272.860 0.000 273.980 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER metal4 ;
  RECT 264.180 0.000 265.300 1.120 ;
  LAYER metal3 ;
  RECT 264.180 0.000 265.300 1.120 ;
  LAYER metal2 ;
  RECT 264.180 0.000 265.300 1.120 ;
  LAYER metal1 ;
  RECT 264.180 0.000 265.300 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER metal4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER metal4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER metal4 ;
  RECT 216.440 0.000 217.560 1.120 ;
  LAYER metal3 ;
  RECT 216.440 0.000 217.560 1.120 ;
  LAYER metal2 ;
  RECT 216.440 0.000 217.560 1.120 ;
  LAYER metal1 ;
  RECT 216.440 0.000 217.560 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER metal4 ;
  RECT 207.760 0.000 208.880 1.120 ;
  LAYER metal3 ;
  RECT 207.760 0.000 208.880 1.120 ;
  LAYER metal2 ;
  RECT 207.760 0.000 208.880 1.120 ;
  LAYER metal1 ;
  RECT 207.760 0.000 208.880 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER metal4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER metal4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI4
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 189.160 0.000 190.280 1.120 ;
  LAYER metal3 ;
  RECT 189.160 0.000 190.280 1.120 ;
  LAYER metal2 ;
  RECT 189.160 0.000 190.280 1.120 ;
  LAYER metal1 ;
  RECT 189.160 0.000 190.280 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal3 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal2 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal1 ;
  RECT 187.300 0.000 188.420 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 182.340 0.000 183.460 1.120 ;
  LAYER metal3 ;
  RECT 182.340 0.000 183.460 1.120 ;
  LAYER metal2 ;
  RECT 182.340 0.000 183.460 1.120 ;
  LAYER metal1 ;
  RECT 182.340 0.000 183.460 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER metal4 ;
  RECT 180.480 0.000 181.600 1.120 ;
  LAYER metal3 ;
  RECT 180.480 0.000 181.600 1.120 ;
  LAYER metal2 ;
  RECT 180.480 0.000 181.600 1.120 ;
  LAYER metal1 ;
  RECT 180.480 0.000 181.600 1.120 ;
 END
END CS
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 178.620 0.000 179.740 1.120 ;
  LAYER metal3 ;
  RECT 178.620 0.000 179.740 1.120 ;
  LAYER metal2 ;
  RECT 178.620 0.000 179.740 1.120 ;
  LAYER metal1 ;
  RECT 178.620 0.000 179.740 1.120 ;
 END
END A3
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 158.780 0.000 159.900 1.120 ;
  LAYER metal3 ;
  RECT 158.780 0.000 159.900 1.120 ;
  LAYER metal2 ;
  RECT 158.780 0.000 159.900 1.120 ;
  LAYER metal1 ;
  RECT 158.780 0.000 159.900 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER metal4 ;
  RECT 155.680 0.000 156.800 1.120 ;
  LAYER metal3 ;
  RECT 155.680 0.000 156.800 1.120 ;
  LAYER metal2 ;
  RECT 155.680 0.000 156.800 1.120 ;
  LAYER metal1 ;
  RECT 155.680 0.000 156.800 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 153.200 0.000 154.320 1.120 ;
  LAYER metal3 ;
  RECT 153.200 0.000 154.320 1.120 ;
  LAYER metal2 ;
  RECT 153.200 0.000 154.320 1.120 ;
  LAYER metal1 ;
  RECT 153.200 0.000 154.320 1.120 ;
 END
END A0
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER metal3 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER metal2 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER metal1 ;
  RECT 148.860 0.000 149.980 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER metal3 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER metal2 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER metal1 ;
  RECT 141.420 0.000 142.540 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER metal3 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER metal2 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER metal1 ;
  RECT 138.320 0.000 139.440 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER metal3 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER metal2 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER metal1 ;
  RECT 130.880 0.000 132.000 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 127.780 0.000 128.900 1.120 ;
  LAYER metal3 ;
  RECT 127.780 0.000 128.900 1.120 ;
  LAYER metal2 ;
  RECT 127.780 0.000 128.900 1.120 ;
  LAYER metal1 ;
  RECT 127.780 0.000 128.900 1.120 ;
 END
END A8
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER metal4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER metal4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER metal4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER metal4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER metal4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER metal4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.059 ;
 PORT
  LAYER metal4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.021 ;
 PORT
  LAYER metal4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 316.200 201.040 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 316.200 201.040 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 316.200 201.040 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 316.200 201.040 ;
  LAYER via ;
  RECT 0.000 0.140 316.200 201.040 ;
  LAYER via2 ;
  RECT 0.000 0.140 316.200 201.040 ;
  LAYER via3 ;
  RECT 0.000 0.140 316.200 201.040 ;
END
END MEM5x5
END LIBRARY



